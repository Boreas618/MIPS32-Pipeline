module Core (
    input clk,
    input rst,
    output write_enabled,
    input [31:0] r_data,
    output [31:0] addr,
    output [31:0] w_data
);

endmodule
